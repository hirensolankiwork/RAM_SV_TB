
package ram_package;

  `include "ram_transaction.sv"
  `include "ram_generator.sv"
  `include "ram_driver.sv"
  `include "ram_monitor.sv"
  `include "ram_env.sv"
  `include "ram_test.sv"

endpackage
